package MergeFifo

module MergeFifo;
endmodule

endpackage : MergeFifo