package Crossbar;

module mkCrossbar #()();

endmodule

endpackage : Crossbar