package TilelinkTracker;



module mkTilelinkTracker();

endmodule

endpackage